LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LUT_mul2 IS
    PORT (
        byte_in : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        byte_out : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END LUT_mul2;

ARCHITECTURE Behavioral OF LUT_mul2 IS
BEGIN
    PROCESS (byte_in) IS
    BEGIN
        CASE byte_in IS
            WHEN x"00" => byte_out <= x"00";
            WHEN x"01" => byte_out <= x"02";
            WHEN x"02" => byte_out <= x"04";
            WHEN x"03" => byte_out <= x"06";
            WHEN x"04" => byte_out <= x"08";
            WHEN x"05" => byte_out <= x"0a";
            WHEN x"06" => byte_out <= x"0c";
            WHEN x"07" => byte_out <= x"0e";
            WHEN x"08" => byte_out <= x"10";
            WHEN x"09" => byte_out <= x"12";
            WHEN x"0a" => byte_out <= x"14";
            WHEN x"0b" => byte_out <= x"16";
            WHEN x"0c" => byte_out <= x"18";
            WHEN x"0d" => byte_out <= x"1a";
            WHEN x"0e" => byte_out <= x"1c";
            WHEN x"0f" => byte_out <= x"1e";
            WHEN x"10" => byte_out <= x"20";
            WHEN x"11" => byte_out <= x"22";
            WHEN x"12" => byte_out <= x"24";
            WHEN x"13" => byte_out <= x"26";
            WHEN x"14" => byte_out <= x"28";
            WHEN x"15" => byte_out <= x"2a";
            WHEN x"16" => byte_out <= x"2c";
            WHEN x"17" => byte_out <= x"2e";
            WHEN x"18" => byte_out <= x"30";
            WHEN x"19" => byte_out <= x"32";
            WHEN x"1a" => byte_out <= x"34";
            WHEN x"1b" => byte_out <= x"36";
            WHEN x"1c" => byte_out <= x"38";
            WHEN x"1d" => byte_out <= x"3a";
            WHEN x"1e" => byte_out <= x"3c";
            WHEN x"1f" => byte_out <= x"3e";
            WHEN x"20" => byte_out <= x"40";
            WHEN x"21" => byte_out <= x"42";
            WHEN x"22" => byte_out <= x"44";
            WHEN x"23" => byte_out <= x"46";
            WHEN x"24" => byte_out <= x"48";
            WHEN x"25" => byte_out <= x"4a";
            WHEN x"26" => byte_out <= x"4c";
            WHEN x"27" => byte_out <= x"4e";
            WHEN x"28" => byte_out <= x"50";
            WHEN x"29" => byte_out <= x"52";
            WHEN x"2a" => byte_out <= x"54";
            WHEN x"2b" => byte_out <= x"56";
            WHEN x"2c" => byte_out <= x"58";
            WHEN x"2d" => byte_out <= x"5a";
            WHEN x"2e" => byte_out <= x"5c";
            WHEN x"2f" => byte_out <= x"5e";
            WHEN x"30" => byte_out <= x"60";
            WHEN x"31" => byte_out <= x"62";
            WHEN x"32" => byte_out <= x"64";
            WHEN x"33" => byte_out <= x"66";
            WHEN x"34" => byte_out <= x"68";
            WHEN x"35" => byte_out <= x"6a";
            WHEN x"36" => byte_out <= x"6c";
            WHEN x"37" => byte_out <= x"6e";
            WHEN x"38" => byte_out <= x"70";
            WHEN x"39" => byte_out <= x"72";
            WHEN x"3a" => byte_out <= x"74";
            WHEN x"3b" => byte_out <= x"76";
            WHEN x"3c" => byte_out <= x"78";
            WHEN x"3d" => byte_out <= x"7a";
            WHEN x"3e" => byte_out <= x"7c";
            WHEN x"3f" => byte_out <= x"7e";
            WHEN x"40" => byte_out <= x"80";
            WHEN x"41" => byte_out <= x"82";
            WHEN x"42" => byte_out <= x"84";
            WHEN x"43" => byte_out <= x"86";
            WHEN x"44" => byte_out <= x"88";
            WHEN x"45" => byte_out <= x"8a";
            WHEN x"46" => byte_out <= x"8c";
            WHEN x"47" => byte_out <= x"8e";
            WHEN x"48" => byte_out <= x"90";
            WHEN x"49" => byte_out <= x"92";
            WHEN x"4a" => byte_out <= x"94";
            WHEN x"4b" => byte_out <= x"96";
            WHEN x"4c" => byte_out <= x"98";
            WHEN x"4d" => byte_out <= x"9a";
            WHEN x"4e" => byte_out <= x"9c";
            WHEN x"4f" => byte_out <= x"9e";
            WHEN x"50" => byte_out <= x"a0";
            WHEN x"51" => byte_out <= x"a2";
            WHEN x"52" => byte_out <= x"a4";
            WHEN x"53" => byte_out <= x"a6";
            WHEN x"54" => byte_out <= x"a8";
            WHEN x"55" => byte_out <= x"aa";
            WHEN x"56" => byte_out <= x"ac";
            WHEN x"57" => byte_out <= x"ae";
            WHEN x"58" => byte_out <= x"b0";
            WHEN x"59" => byte_out <= x"b2";
            WHEN x"5a" => byte_out <= x"b4";
            WHEN x"5b" => byte_out <= x"b6";
            WHEN x"5c" => byte_out <= x"b8";
            WHEN x"5d" => byte_out <= x"ba";
            WHEN x"5e" => byte_out <= x"bc";
            WHEN x"5f" => byte_out <= x"be";
            WHEN x"60" => byte_out <= x"c0";
            WHEN x"61" => byte_out <= x"c2";
            WHEN x"62" => byte_out <= x"c4";
            WHEN x"63" => byte_out <= x"c6";
            WHEN x"64" => byte_out <= x"c8";
            WHEN x"65" => byte_out <= x"ca";
            WHEN x"66" => byte_out <= x"cc";
            WHEN x"67" => byte_out <= x"ce";
            WHEN x"68" => byte_out <= x"d0";
            WHEN x"69" => byte_out <= x"d2";
            WHEN x"6a" => byte_out <= x"d4";
            WHEN x"6b" => byte_out <= x"d6";
            WHEN x"6c" => byte_out <= x"d8";
            WHEN x"6d" => byte_out <= x"da";
            WHEN x"6e" => byte_out <= x"dc";
            WHEN x"6f" => byte_out <= x"de";
            WHEN x"70" => byte_out <= x"e0";
            WHEN x"71" => byte_out <= x"e2";
            WHEN x"72" => byte_out <= x"e4";
            WHEN x"73" => byte_out <= x"e6";
            WHEN x"74" => byte_out <= x"e8";
            WHEN x"75" => byte_out <= x"ea";
            WHEN x"76" => byte_out <= x"ec";
            WHEN x"77" => byte_out <= x"ee";
            WHEN x"78" => byte_out <= x"f0";
            WHEN x"79" => byte_out <= x"f2";
            WHEN x"7a" => byte_out <= x"f4";
            WHEN x"7b" => byte_out <= x"f6";
            WHEN x"7c" => byte_out <= x"f8";
            WHEN x"7d" => byte_out <= x"fa";
            WHEN x"7e" => byte_out <= x"fc";
            WHEN x"7f" => byte_out <= x"fe";
            WHEN x"80" => byte_out <= x"1b";
            WHEN x"81" => byte_out <= x"19";
            WHEN x"82" => byte_out <= x"1f";
            WHEN x"83" => byte_out <= x"1d";
            WHEN x"84" => byte_out <= x"13";
            WHEN x"85" => byte_out <= x"11";
            WHEN x"86" => byte_out <= x"17";
            WHEN x"87" => byte_out <= x"15";
            WHEN x"88" => byte_out <= x"0b";
            WHEN x"89" => byte_out <= x"09";
            WHEN x"8a" => byte_out <= x"0f";
            WHEN x"8b" => byte_out <= x"0d";
            WHEN x"8c" => byte_out <= x"03";
            WHEN x"8d" => byte_out <= x"01";
            WHEN x"8e" => byte_out <= x"07";
            WHEN x"8f" => byte_out <= x"05";
            WHEN x"90" => byte_out <= x"3b";
            WHEN x"91" => byte_out <= x"39";
            WHEN x"92" => byte_out <= x"3f";
            WHEN x"93" => byte_out <= x"3d";
            WHEN x"94" => byte_out <= x"33";
            WHEN x"95" => byte_out <= x"31";
            WHEN x"96" => byte_out <= x"37";
            WHEN x"97" => byte_out <= x"35";
            WHEN x"98" => byte_out <= x"2b";
            WHEN x"99" => byte_out <= x"29";
            WHEN x"9a" => byte_out <= x"2f";
            WHEN x"9b" => byte_out <= x"2d";
            WHEN x"9c" => byte_out <= x"23";
            WHEN x"9d" => byte_out <= x"21";
            WHEN x"9e" => byte_out <= x"27";
            WHEN x"9f" => byte_out <= x"25";
            WHEN x"a0" => byte_out <= x"5b";
            WHEN x"a1" => byte_out <= x"59";
            WHEN x"a2" => byte_out <= x"5f";
            WHEN x"a3" => byte_out <= x"5d";
            WHEN x"a4" => byte_out <= x"53";
            WHEN x"a5" => byte_out <= x"51";
            WHEN x"a6" => byte_out <= x"57";
            WHEN x"a7" => byte_out <= x"55";
            WHEN x"a8" => byte_out <= x"4b";
            WHEN x"a9" => byte_out <= x"49";
            WHEN x"aa" => byte_out <= x"4f";
            WHEN x"ab" => byte_out <= x"4d";
            WHEN x"ac" => byte_out <= x"43";
            WHEN x"ad" => byte_out <= x"41";
            WHEN x"ae" => byte_out <= x"47";
            WHEN x"af" => byte_out <= x"45";
            WHEN x"b0" => byte_out <= x"7b";
            WHEN x"b1" => byte_out <= x"79";
            WHEN x"b2" => byte_out <= x"7f";
            WHEN x"b3" => byte_out <= x"7d";
            WHEN x"b4" => byte_out <= x"73";
            WHEN x"b5" => byte_out <= x"71";
            WHEN x"b6" => byte_out <= x"77";
            WHEN x"b7" => byte_out <= x"75";
            WHEN x"b8" => byte_out <= x"6b";
            WHEN x"b9" => byte_out <= x"69";
            WHEN x"ba" => byte_out <= x"6f";
            WHEN x"bb" => byte_out <= x"6d";
            WHEN x"bc" => byte_out <= x"63";
            WHEN x"bd" => byte_out <= x"61";
            WHEN x"be" => byte_out <= x"67";
            WHEN x"bf" => byte_out <= x"65";
            WHEN x"c0" => byte_out <= x"9b";
            WHEN x"c1" => byte_out <= x"99";
            WHEN x"c2" => byte_out <= x"9f";
            WHEN x"c3" => byte_out <= x"9d";
            WHEN x"c4" => byte_out <= x"93";
            WHEN x"c5" => byte_out <= x"91";
            WHEN x"c6" => byte_out <= x"97";
            WHEN x"c7" => byte_out <= x"95";
            WHEN x"c8" => byte_out <= x"8b";
            WHEN x"c9" => byte_out <= x"89";
            WHEN x"ca" => byte_out <= x"8f";
            WHEN x"cb" => byte_out <= x"8d";
            WHEN x"cc" => byte_out <= x"83";
            WHEN x"cd" => byte_out <= x"81";
            WHEN x"ce" => byte_out <= x"87";
            WHEN x"cf" => byte_out <= x"85";
            WHEN x"d0" => byte_out <= x"bb";
            WHEN x"d1" => byte_out <= x"b9";
            WHEN x"d2" => byte_out <= x"bf";
            WHEN x"d3" => byte_out <= x"bd";
            WHEN x"d4" => byte_out <= x"b3";
            WHEN x"d5" => byte_out <= x"b1";
            WHEN x"d6" => byte_out <= x"b7";
            WHEN x"d7" => byte_out <= x"b5";
            WHEN x"d8" => byte_out <= x"ab";
            WHEN x"d9" => byte_out <= x"a9";
            WHEN x"da" => byte_out <= x"af";
            WHEN x"db" => byte_out <= x"ad";
            WHEN x"dc" => byte_out <= x"a3";
            WHEN x"dd" => byte_out <= x"a1";
            WHEN x"de" => byte_out <= x"a7";
            WHEN x"df" => byte_out <= x"a5";
            WHEN x"e0" => byte_out <= x"db";
            WHEN x"e1" => byte_out <= x"d9";
            WHEN x"e2" => byte_out <= x"df";
            WHEN x"e3" => byte_out <= x"dd";
            WHEN x"e4" => byte_out <= x"d3";
            WHEN x"e5" => byte_out <= x"d1";
            WHEN x"e6" => byte_out <= x"d7";
            WHEN x"e7" => byte_out <= x"d5";
            WHEN x"e8" => byte_out <= x"cb";
            WHEN x"e9" => byte_out <= x"c9";
            WHEN x"ea" => byte_out <= x"cf";
            WHEN x"eb" => byte_out <= x"cd";
            WHEN x"ec" => byte_out <= x"c3";
            WHEN x"ed" => byte_out <= x"c1";
            WHEN x"ee" => byte_out <= x"c7";
            WHEN x"ef" => byte_out <= x"c5";
            WHEN x"f0" => byte_out <= x"fb";
            WHEN x"f1" => byte_out <= x"f9";
            WHEN x"f2" => byte_out <= x"ff";
            WHEN x"f3" => byte_out <= x"fd";
            WHEN x"f4" => byte_out <= x"f3";
            WHEN x"f5" => byte_out <= x"f1";
            WHEN x"f6" => byte_out <= x"f7";
            WHEN x"f7" => byte_out <= x"f5";
            WHEN x"f8" => byte_out <= x"eb";
            WHEN x"f9" => byte_out <= x"e9";
            WHEN x"fa" => byte_out <= x"ef";
            WHEN x"fb" => byte_out <= x"ed";
            WHEN x"fc" => byte_out <= x"e3";
            WHEN x"fd" => byte_out <= x"e1";
            WHEN x"fe" => byte_out <= x"e7";
            WHEN x"ff" => byte_out <= x"e5";
            WHEN OTHERS => byte_out <= x"00";
        END CASE;
    END PROCESS;

END Behavioral;