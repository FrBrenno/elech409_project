library ieee;
use ieee.std_logic_1164.all;

entity AES_encryption_tb is
end AES_encryption_tb;

architecture tb_arch of AES_encryption_tb is

begin

end tb_arch;
